module Adder (
    input  signed [37:0] in1,
    in2,
    output signed [37:0] out
);
  assign out = in1 + in2;
endmodule

